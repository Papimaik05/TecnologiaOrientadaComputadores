    Mac OS X            	   2   �      �                                      ATTR       �   �   3                  �     com.apple.lastuseddate#PS       �   #  com.apple.quarantine }_�a    !O8    q/0082;61a35d06;The\x20Unarchiver; 