    Mac OS X            	   2  {     �                                      ATTR      �   �   �                  �   �  "com.apple.LaunchServices.OpenWith      z     com.apple.lastuseddate#PS      �   #  com.apple.quarantine bplist00�WversionTpath_bundleidentifier _/Applications/BBEdit.app_com.barebones.bbedit/1L                            c�_�a    $y�    q/00e2;61a35d06;The\x20Unarchiver; 